module testbench();
	logic        clk, reset;
	logic        n, s, e, w, win, die, winexpected, dieexpected;
	logic [31:0] vectornum, errors;
	logic [5:0]  testvectors[10000:0];
	
	// задание (определение) тестируемого устройства
	game dut(clk, reset, n, s, e, w, win, die); 

	// Тактовый генератор
	always
		begin
			clk=1; #5; 
			clk=0; #5; 
		end
	
	// при старте теста загрузить векторы и дать импульс сброса
	initial 
		begin
			$readmemb("game.tv", testvectors); 
			vectornum = 0; 
			errors = 0;
			reset = 1; #22; 
			reset = 0; #70;
			reset = 1; #10;
			reset = 0; #70;
			reset = 1; #10;
			reset = 0;
		end 
		
	// подать тестовые векторы по переднему(нарстающему) фронту такта
	always @(posedge clk) 
		begin
			#1; 
			{n, s, e, w, winexpected, dieexpected} = testvectors[vectornum]; 
		end 
	
	// проверить результаты по заднему(спадающему) фронту такта
	always @(negedge clk) 
		if (~reset) 
			begin    // пропустить проверку при сбросе
				if (win !== winexpected || die !== dieexpected) 
					begin // проверить результаты
						$display("Error: inputs = %b", {n, s, e, w});
						$display(" outputs = %b %b (%b %b expected)", 
							win, die, winexpected, dieexpected); 
						errors = errors + 1; 
					end

				vectornum = vectornum + 1;
				if (testvectors[vectornum] === 6'bx) 
					begin 
						$display("%d tests completed with %d errors", vectornum, errors); 
						$stop; 
					end 
			end 
	
endmodule 