// Поведенческий Verilog объясняет взаимоотношения между вводами и выводами
// К примеру: assign y = a & b;
// Структурный Verilog описывает структуры сформированные более простыми компонентами
// К примеру: and g1(y, a, b);
// Разделы 4.1-4.3 в книге (начиная со стр. 171) описывают эти 
// различия в деталях

// Этот модуль структурный или поведенческий?
module fulladder(input  logic a, b, cin,
		     output logic sum, cout);
	
	// Объявить 5 внутренних логических сигналов или локальных переменных, 
	// которые могут использоваться только в пределах этого модуля
	logic ns, n1, n2, n3, n4;
	
	// Следующие логические вентили являются частью спецификации SystemVerilog
	// (встроенные примитивы).
	// Первый сигнал (к примеру, ns) является выводом. Остальные(e.g., a, b) являются 
	// вводами.

	// sum logic
	xor x1(ns, a, b);		// ns = a XOR b
	xor x2(sum, ns, cin);	// sum = ns XOR cin
	
	// carry logic
	and a1(n1, a, b);		// n1 = a & b
	and a2(n2, a, cin);		// n2 = a & cin
	and a3(n3, b, cin);		// n3 = b & cin
	or o1(n4, n1, n2);		// n4 = n1 | n2
	or o2(cout, n3, n4);	// cout = n3 | n4

// Этот пример является структурным Verilog'ом, поскольку модуль описан 
// структурно, используя более фундаментальные блоки построения 
endmodule